`timescale 1ns/1ns
module Shifter( dataA, dataB, dataOut, reset);
  input reset;
  input [31:0] dataA;
  input [31:0] dataB;
  output [31:0] dataOut;

  wire [31:0] SHAMT1, SHAMT2, SHAMT3, SHAMT4;
  wire [31:0] temp;

  wire reset_wire;

  // Level 1
  MUX2_1 mux0( .i0(dataA[0]), .i1(dataA[1]), .sel(dataB[0]), .out(SHAMT1[0]) ) ;
  MUX2_1 mux1( .i0(dataA[1]), .i1(dataA[2]), .sel(dataB[0]), .out(SHAMT1[1]) ) ;
  MUX2_1 mux2( .i0(dataA[2]), .i1(dataA[3]), .sel(dataB[0]), .out(SHAMT1[2]) ) ;
  MUX2_1 mux3( .i0(dataA[3]), .i1(dataA[4]), .sel(dataB[0]), .out(SHAMT1[3]) ) ;
  MUX2_1 mux4( .i0(dataA[4]), .i1(dataA[5]), .sel(dataB[0]), .out(SHAMT1[4]) ) ;
  MUX2_1 mux5( .i0(dataA[5]), .i1(dataA[6]), .sel(dataB[0]), .out(SHAMT1[5]) ) ;
  MUX2_1 mux6( .i0(dataA[6]), .i1(dataA[7]), .sel(dataB[0]), .out(SHAMT1[6]) ) ;
  MUX2_1 mux7( .i0(dataA[7]), .i1(dataA[8]), .sel(dataB[0]), .out(SHAMT1[7]) ) ;
  MUX2_1 mux8( .i0(dataA[8]), .i1(dataA[9]), .sel(dataB[0]), .out(SHAMT1[8]) ) ;
  MUX2_1 mux9( .i0(dataA[9]), .i1(dataA[10]), .sel(dataB[0]), .out(SHAMT1[9]) ) ;
  MUX2_1 mux10( .i0(dataA[10]), .i1(dataA[11]), .sel(dataB[0]), .out(SHAMT1[10]) ) ;
  MUX2_1 mux11( .i0(dataA[11]), .i1(dataA[12]), .sel(dataB[0]), .out(SHAMT1[11]) ) ;
  MUX2_1 mux12( .i0(dataA[12]), .i1(dataA[13]), .sel(dataB[0]), .out(SHAMT1[12]) ) ;
  MUX2_1 mux13( .i0(dataA[13]), .i1(dataA[14]), .sel(dataB[0]), .out(SHAMT1[13]) ) ;
  MUX2_1 mux14( .i0(dataA[14]), .i1(dataA[15]), .sel(dataB[0]), .out(SHAMT1[14]) ) ;
  MUX2_1 mux15( .i0(dataA[15]), .i1(dataA[16]), .sel(dataB[0]), .out(SHAMT1[15]) ) ;
  MUX2_1 mux16( .i0(dataA[16]), .i1(dataA[17]), .sel(dataB[0]), .out(SHAMT1[16]) ) ;
  MUX2_1 mux17( .i0(dataA[17]), .i1(dataA[18]), .sel(dataB[0]), .out(SHAMT1[17]) ) ;
  MUX2_1 mux18( .i0(dataA[18]), .i1(dataA[19]), .sel(dataB[0]), .out(SHAMT1[18]) ) ;
  MUX2_1 mux19( .i0(dataA[19]), .i1(dataA[20]), .sel(dataB[0]), .out(SHAMT1[19]) ) ;
  MUX2_1 mux20( .i0(dataA[20]), .i1(dataA[21]), .sel(dataB[0]), .out(SHAMT1[20]) ) ;
  MUX2_1 mux21( .i0(dataA[21]), .i1(dataA[22]), .sel(dataB[0]), .out(SHAMT1[21]) ) ;
  MUX2_1 mux22( .i0(dataA[22]), .i1(dataA[23]), .sel(dataB[0]), .out(SHAMT1[22]) ) ;
  MUX2_1 mux23( .i0(dataA[23]), .i1(dataA[24]), .sel(dataB[0]), .out(SHAMT1[23]) ) ;
  MUX2_1 mux24( .i0(dataA[24]), .i1(dataA[25]), .sel(dataB[0]), .out(SHAMT1[24]) ) ;
  MUX2_1 mux25( .i0(dataA[25]), .i1(dataA[26]), .sel(dataB[0]), .out(SHAMT1[25]) ) ;
  MUX2_1 mux26( .i0(dataA[26]), .i1(dataA[27]), .sel(dataB[0]), .out(SHAMT1[26]) ) ;
  MUX2_1 mux27( .i0(dataA[27]), .i1(dataA[28]), .sel(dataB[0]), .out(SHAMT1[27]) ) ;
  MUX2_1 mux28( .i0(dataA[28]), .i1(dataA[29]), .sel(dataB[0]), .out(SHAMT1[28]) ) ;
  MUX2_1 mux29( .i0(dataA[29]), .i1(dataA[30]), .sel(dataB[0]), .out(SHAMT1[29]) ) ;
  MUX2_1 mux30( .i0(dataA[30]), .i1(dataA[31]), .sel(dataB[0]), .out(SHAMT1[30]) ) ;
  MUX2_1 mux31( .i0(dataA[31]), .i1(1'b0), .sel(dataB[0]), .out(SHAMT1[31]) ) ;

  // Level 2
  MUX2_1 mux00( .i0(SHAMT1[0]), .i1(SHAMT1[2]), .sel(dataB[1]), .out(SHAMT2[0]) ) ;
  MUX2_1 mux01( .i0(SHAMT1[1]), .i1(SHAMT1[3]), .sel(dataB[1]), .out(SHAMT2[1]) ) ;
  MUX2_1 mux02( .i0(SHAMT1[2]), .i1(SHAMT1[4]), .sel(dataB[1]), .out(SHAMT2[2]) ) ;
  MUX2_1 mux03( .i0(SHAMT1[3]), .i1(SHAMT1[5]), .sel(dataB[1]), .out(SHAMT2[3]) ) ;
  MUX2_1 mux04( .i0(SHAMT1[4]), .i1(SHAMT1[6]), .sel(dataB[1]), .out(SHAMT2[4]) ) ;
  MUX2_1 mux05( .i0(SHAMT1[5]), .i1(SHAMT1[7]), .sel(dataB[1]), .out(SHAMT2[5]) ) ;
  MUX2_1 mux06( .i0(SHAMT1[6]), .i1(SHAMT1[8]), .sel(dataB[1]), .out(SHAMT2[6]) ) ;
  MUX2_1 mux07( .i0(SHAMT1[7]), .i1(SHAMT1[9]), .sel(dataB[1]), .out(SHAMT2[7]) ) ;
  MUX2_1 mux08( .i0(SHAMT1[8]), .i1(SHAMT1[10]), .sel(dataB[1]), .out(SHAMT2[8]) ) ;
  MUX2_1 mux09( .i0(SHAMT1[9]), .i1(SHAMT1[11]), .sel(dataB[1]), .out(SHAMT2[9]) ) ;
  MUX2_1 mux010( .i0(SHAMT1[10]), .i1(SHAMT1[12]), .sel(dataB[1]), .out(SHAMT2[10]) ) ;
  MUX2_1 mux011( .i0(SHAMT1[11]), .i1(SHAMT1[13]), .sel(dataB[1]), .out(SHAMT2[11]) ) ;
  MUX2_1 mux012( .i0(SHAMT1[12]), .i1(SHAMT1[14]), .sel(dataB[1]), .out(SHAMT2[12]) ) ;
  MUX2_1 mux013( .i0(SHAMT1[13]), .i1(SHAMT1[15]), .sel(dataB[1]), .out(SHAMT2[13]) ) ;
  MUX2_1 mux014( .i0(SHAMT1[14]), .i1(SHAMT1[16]), .sel(dataB[1]), .out(SHAMT2[14]) ) ;
  MUX2_1 mux015( .i0(SHAMT1[15]), .i1(SHAMT1[17]), .sel(dataB[1]), .out(SHAMT2[15]) ) ;
  MUX2_1 mux016( .i0(SHAMT1[16]), .i1(SHAMT1[18]), .sel(dataB[1]), .out(SHAMT2[16]) ) ;
  MUX2_1 mux017( .i0(SHAMT1[17]), .i1(SHAMT1[19]), .sel(dataB[1]), .out(SHAMT2[17]) ) ;
  MUX2_1 mux018( .i0(SHAMT1[18]), .i1(SHAMT1[20]), .sel(dataB[1]), .out(SHAMT2[18]) ) ;
  MUX2_1 mux019( .i0(SHAMT1[19]), .i1(SHAMT1[21]), .sel(dataB[1]), .out(SHAMT2[19]) ) ;
  MUX2_1 mux020( .i0(SHAMT1[20]), .i1(SHAMT1[22]), .sel(dataB[1]), .out(SHAMT2[20]) ) ;
  MUX2_1 mux021( .i0(SHAMT1[21]), .i1(SHAMT1[23]), .sel(dataB[1]), .out(SHAMT2[21]) ) ;
  MUX2_1 mux022( .i0(SHAMT1[22]), .i1(SHAMT1[24]), .sel(dataB[1]), .out(SHAMT2[22]) ) ;
  MUX2_1 mux023( .i0(SHAMT1[23]), .i1(SHAMT1[25]), .sel(dataB[1]), .out(SHAMT2[23]) ) ;
  MUX2_1 mux024( .i0(SHAMT1[24]), .i1(SHAMT1[26]), .sel(dataB[1]), .out(SHAMT2[24]) ) ;
  MUX2_1 mux025( .i0(SHAMT1[25]), .i1(SHAMT1[27]), .sel(dataB[1]), .out(SHAMT2[25]) ) ;
  MUX2_1 mux026( .i0(SHAMT1[26]), .i1(SHAMT1[28]), .sel(dataB[1]), .out(SHAMT2[26]) ) ;
  MUX2_1 mux027( .i0(SHAMT1[27]), .i1(SHAMT1[29]), .sel(dataB[1]), .out(SHAMT2[27]) ) ;
  MUX2_1 mux028( .i0(SHAMT1[28]), .i1(SHAMT1[30]), .sel(dataB[1]), .out(SHAMT2[28]) ) ;
  MUX2_1 mux029( .i0(SHAMT1[29]), .i1(SHAMT1[31]), .sel(dataB[1]), .out(SHAMT2[29]) ) ;
  MUX2_1 mux030( .i0(SHAMT1[30]), .i1(1'b0), .sel(dataB[1]), .out(SHAMT2[30]) ) ;
  MUX2_1 mux031( .i0(SHAMT1[31]), .i1(1'b0), .sel(dataB[1]), .out(SHAMT2[31]) ) ;

  // Level 3
  MUX2_1 mux000( .i0(SHAMT2[0]), .i1(SHAMT2[4]), .sel(dataB[2]), .out(SHAMT3[0]) ) ;
  MUX2_1 mux001( .i0(SHAMT2[1]), .i1(SHAMT2[5]), .sel(dataB[2]), .out(SHAMT3[1]) ) ;
  MUX2_1 mux002( .i0(SHAMT2[2]), .i1(SHAMT2[6]), .sel(dataB[2]), .out(SHAMT3[2]) ) ;
  MUX2_1 mux003( .i0(SHAMT2[3]), .i1(SHAMT2[7]), .sel(dataB[2]), .out(SHAMT3[3]) ) ;
  MUX2_1 mux004( .i0(SHAMT2[4]), .i1(SHAMT2[8]), .sel(dataB[2]), .out(SHAMT3[4]) ) ;
  MUX2_1 mux005( .i0(SHAMT2[5]), .i1(SHAMT2[9]), .sel(dataB[2]), .out(SHAMT3[5]) ) ;
  MUX2_1 mux006( .i0(SHAMT2[6]), .i1(SHAMT2[10]), .sel(dataB[2]), .out(SHAMT3[6]) ) ;
  MUX2_1 mux007( .i0(SHAMT2[7]), .i1(SHAMT2[11]), .sel(dataB[2]), .out(SHAMT3[7]) ) ;
  MUX2_1 mux008( .i0(SHAMT2[8]), .i1(SHAMT2[12]), .sel(dataB[2]), .out(SHAMT3[8]) ) ;
  MUX2_1 mux009( .i0(SHAMT2[9]), .i1(SHAMT2[13]), .sel(dataB[2]), .out(SHAMT3[9]) ) ;
  MUX2_1 mux0010( .i0(SHAMT2[10]), .i1(SHAMT2[14]), .sel(dataB[2]), .out(SHAMT3[10]) ) ;
  MUX2_1 mux0011( .i0(SHAMT2[11]), .i1(SHAMT2[15]), .sel(dataB[2]), .out(SHAMT3[11]) ) ;
  MUX2_1 mux0012( .i0(SHAMT2[12]), .i1(SHAMT2[16]), .sel(dataB[2]), .out(SHAMT3[12]) ) ;
  MUX2_1 mux0013( .i0(SHAMT2[13]), .i1(SHAMT2[17]), .sel(dataB[2]), .out(SHAMT3[13]) ) ;
  MUX2_1 mux0014( .i0(SHAMT2[14]), .i1(SHAMT2[18]), .sel(dataB[2]), .out(SHAMT3[14]) ) ;
  MUX2_1 mux0015( .i0(SHAMT2[15]), .i1(SHAMT2[19]), .sel(dataB[2]), .out(SHAMT3[15]) ) ;
  MUX2_1 mux0016( .i0(SHAMT2[16]), .i1(SHAMT2[20]), .sel(dataB[2]), .out(SHAMT3[16]) ) ;
  MUX2_1 mux0017( .i0(SHAMT2[17]), .i1(SHAMT2[21]), .sel(dataB[2]), .out(SHAMT3[17]) ) ;
  MUX2_1 mux0018( .i0(SHAMT2[18]), .i1(SHAMT2[22]), .sel(dataB[2]), .out(SHAMT3[18]) ) ;
  MUX2_1 mux0019( .i0(SHAMT2[19]), .i1(SHAMT2[23]), .sel(dataB[2]), .out(SHAMT3[19]) ) ;
  MUX2_1 mux0020( .i0(SHAMT2[20]), .i1(SHAMT2[24]), .sel(dataB[2]), .out(SHAMT3[20]) ) ;
  MUX2_1 mux0021( .i0(SHAMT2[21]), .i1(SHAMT2[25]), .sel(dataB[2]), .out(SHAMT3[21]) ) ;
  MUX2_1 mux0022( .i0(SHAMT2[22]), .i1(SHAMT2[26]), .sel(dataB[2]), .out(SHAMT3[22]) ) ;
  MUX2_1 mux0023( .i0(SHAMT2[23]), .i1(SHAMT2[27]), .sel(dataB[2]), .out(SHAMT3[23]) ) ;
  MUX2_1 mux0024( .i0(SHAMT2[24]), .i1(SHAMT2[28]), .sel(dataB[2]), .out(SHAMT3[24]) ) ;
  MUX2_1 mux0025( .i0(SHAMT2[25]), .i1(SHAMT2[29]), .sel(dataB[2]), .out(SHAMT3[25]) ) ;
  MUX2_1 mux0026( .i0(SHAMT2[26]), .i1(SHAMT2[30]), .sel(dataB[2]), .out(SHAMT3[26]) ) ;
  MUX2_1 mux0027( .i0(SHAMT2[27]), .i1(SHAMT2[31]), .sel(dataB[2]), .out(SHAMT3[27]) ) ;
  MUX2_1 mux0028( .i0(SHAMT2[28]), .i1(1'b0), .sel(dataB[2]), .out(SHAMT3[28]) ) ;
  MUX2_1 mux0029( .i0(SHAMT2[29]), .i1(1'b0), .sel(dataB[2]), .out(SHAMT3[29]) ) ;
  MUX2_1 mux0030( .i0(SHAMT2[30]), .i1(1'b0), .sel(dataB[2]), .out(SHAMT3[30]) ) ;
  MUX2_1 mux0031( .i0(SHAMT2[31]), .i1(1'b0), .sel(dataB[2]), .out(SHAMT3[31]) ) ;
        
  // Level 4
  MUX2_1 mux0000( .i0(SHAMT3[0]), .i1(SHAMT3[8]), .sel(dataB[3]), .out(SHAMT4[0]) ) ;
  MUX2_1 mux0001( .i0(SHAMT3[1]), .i1(SHAMT3[9]), .sel(dataB[3]), .out(SHAMT4[1]) ) ;
  MUX2_1 mux0002( .i0(SHAMT3[2]), .i1(SHAMT3[10]), .sel(dataB[3]), .out(SHAMT4[2]) ) ;
  MUX2_1 mux0003( .i0(SHAMT3[3]), .i1(SHAMT3[11]), .sel(dataB[3]), .out(SHAMT4[3]) ) ;
  MUX2_1 mux0004( .i0(SHAMT3[4]), .i1(SHAMT3[12]), .sel(dataB[3]), .out(SHAMT4[4]) ) ;
  MUX2_1 mux0005( .i0(SHAMT3[5]), .i1(SHAMT3[13]), .sel(dataB[3]), .out(SHAMT4[5]) ) ;
  MUX2_1 mux0006( .i0(SHAMT3[6]), .i1(SHAMT3[14]), .sel(dataB[3]), .out(SHAMT4[6]) ) ;
  MUX2_1 mux0007( .i0(SHAMT3[7]), .i1(SHAMT3[15]), .sel(dataB[3]), .out(SHAMT4[7]) ) ;
  MUX2_1 mux0008( .i0(SHAMT3[8]), .i1(SHAMT3[16]), .sel(dataB[3]), .out(SHAMT4[8]) ) ;
  MUX2_1 mux0009( .i0(SHAMT3[9]), .i1(SHAMT3[17]), .sel(dataB[3]), .out(SHAMT4[9]) ) ;
  MUX2_1 mux00010( .i0(SHAMT3[10]), .i1(SHAMT3[18]), .sel(dataB[3]), .out(SHAMT4[10]) ) ;
  MUX2_1 mux00011( .i0(SHAMT3[11]), .i1(SHAMT3[19]), .sel(dataB[3]), .out(SHAMT4[11]) ) ;
  MUX2_1 mux00012( .i0(SHAMT3[12]), .i1(SHAMT3[20]), .sel(dataB[3]), .out(SHAMT4[12]) ) ;
  MUX2_1 mux00013( .i0(SHAMT3[13]), .i1(SHAMT3[21]), .sel(dataB[3]), .out(SHAMT4[13]) ) ;
  MUX2_1 mux00014( .i0(SHAMT3[14]), .i1(SHAMT3[22]), .sel(dataB[3]), .out(SHAMT4[14]) ) ;
  MUX2_1 mux00015( .i0(SHAMT3[15]), .i1(SHAMT3[23]), .sel(dataB[3]), .out(SHAMT4[15]) ) ;
  MUX2_1 mux00016( .i0(SHAMT3[16]), .i1(SHAMT3[24]), .sel(dataB[3]), .out(SHAMT4[16]) ) ;
  MUX2_1 mux00017( .i0(SHAMT3[17]), .i1(SHAMT3[25]), .sel(dataB[3]), .out(SHAMT4[17]) ) ;
  MUX2_1 mux00018( .i0(SHAMT3[18]), .i1(SHAMT3[26]), .sel(dataB[3]), .out(SHAMT4[18]) ) ;
  MUX2_1 mux00019( .i0(SHAMT3[19]), .i1(SHAMT3[27]), .sel(dataB[3]), .out(SHAMT4[19]) ) ;
  MUX2_1 mux00020( .i0(SHAMT3[20]), .i1(SHAMT3[28]), .sel(dataB[3]), .out(SHAMT4[20]) ) ;
  MUX2_1 mux00021( .i0(SHAMT3[21]), .i1(SHAMT3[29]), .sel(dataB[3]), .out(SHAMT4[21]) ) ;
  MUX2_1 mux00022( .i0(SHAMT3[22]), .i1(SHAMT3[30]), .sel(dataB[3]), .out(SHAMT4[22]) ) ;
  MUX2_1 mux00023( .i0(SHAMT3[23]), .i1(SHAMT3[31]), .sel(dataB[3]), .out(SHAMT4[23]) ) ;
  MUX2_1 mux00024( .i0(SHAMT3[24]), .i1(1'b0), .sel(dataB[3]), .out(SHAMT4[24]) ) ;
  MUX2_1 mux00025( .i0(SHAMT3[25]), .i1(1'b0), .sel(dataB[3]), .out(SHAMT4[25]) ) ;
  MUX2_1 mux00026( .i0(SHAMT3[26]), .i1(1'b0), .sel(dataB[3]), .out(SHAMT4[26]) ) ;
  MUX2_1 mux00027( .i0(SHAMT3[27]), .i1(1'b0), .sel(dataB[3]), .out(SHAMT4[27]) ) ;
  MUX2_1 mux00028( .i0(SHAMT3[28]), .i1(1'b0), .sel(dataB[3]), .out(SHAMT4[28]) ) ;
  MUX2_1 mux00029( .i0(SHAMT3[29]), .i1(1'b0), .sel(dataB[3]), .out(SHAMT4[29]) ) ;
  MUX2_1 mux00030( .i0(SHAMT3[30]), .i1(1'b0), .sel(dataB[3]), .out(SHAMT4[30]) ) ;
  MUX2_1 mux00031( .i0(SHAMT3[31]), .i1(1'b0), .sel(dataB[3]), .out(SHAMT4[31]) ) ;

  // Level 5
  MUX2_1 mux00000( .i0(SHAMT4[0]), .i1(SHAMT4[17]), .sel(dataB[4]), .out(temp[0]) ) ;
  MUX2_1 mux00001( .i0(SHAMT4[1]), .i1(SHAMT4[18]), .sel(dataB[4]), .out(temp[1]) ) ;
  MUX2_1 mux00002( .i0(SHAMT4[2]), .i1(SHAMT4[19]), .sel(dataB[4]), .out(temp[2]) ) ;
  MUX2_1 mux00003( .i0(SHAMT4[3]), .i1(SHAMT4[20]), .sel(dataB[4]), .out(temp[3]) ) ;
  MUX2_1 mux00004( .i0(SHAMT4[4]), .i1(SHAMT4[21]), .sel(dataB[4]), .out(temp[4]) ) ;
  MUX2_1 mux00005( .i0(SHAMT4[5]), .i1(SHAMT4[22]), .sel(dataB[4]), .out(temp[5]) ) ;
  MUX2_1 mux00006( .i0(SHAMT4[6]), .i1(SHAMT4[23]), .sel(dataB[4]), .out(temp[6]) ) ;
  MUX2_1 mux00007( .i0(SHAMT4[7]), .i1(SHAMT4[24]), .sel(dataB[4]), .out(temp[7]) ) ;
  MUX2_1 mux00008( .i0(SHAMT4[8]), .i1(SHAMT4[25]), .sel(dataB[4]), .out(temp[8]) ) ;
  MUX2_1 mux00009( .i0(SHAMT4[9]), .i1(SHAMT4[26]), .sel(dataB[4]), .out(temp[9]) ) ;
  MUX2_1 mux000010( .i0(SHAMT4[10]), .i1(SHAMT4[27]), .sel(dataB[4]), .out(temp[10]) ) ;
  MUX2_1 mux000011( .i0(SHAMT4[11]), .i1(SHAMT4[28]), .sel(dataB[4]), .out(temp[11]) ) ;
  MUX2_1 mux000012( .i0(SHAMT4[12]), .i1(SHAMT4[29]), .sel(dataB[4]), .out(temp[12]) ) ;
  MUX2_1 mux000013( .i0(SHAMT4[13]), .i1(SHAMT4[30]), .sel(dataB[4]), .out(temp[13]) ) ;
  MUX2_1 mux000014( .i0(SHAMT4[14]), .i1(SHAMT4[31]), .sel(dataB[4]), .out(temp[14]) ) ;
  MUX2_1 mux000015( .i0(SHAMT4[15]), .i1(1'b0), .sel(dataB[4]), .out(temp[15]) ) ;
  MUX2_1 mux000016( .i0(SHAMT4[16]), .i1(1'b0), .sel(dataB[4]), .out(temp[16]) ) ;
  MUX2_1 mux000017( .i0(SHAMT4[17]), .i1(1'b0), .sel(dataB[4]), .out(temp[17]) ) ;
  MUX2_1 mux000018( .i0(SHAMT4[18]), .i1(1'b0), .sel(dataB[4]), .out(temp[18]) ) ;
  MUX2_1 mux000019( .i0(SHAMT4[19]), .i1(1'b0), .sel(dataB[4]), .out(temp[19]) ) ;
  MUX2_1 mux000020( .i0(SHAMT4[20]), .i1(1'b0), .sel(dataB[4]), .out(temp[20]) ) ;
  MUX2_1 mux000021( .i0(SHAMT4[21]), .i1(1'b0), .sel(dataB[4]), .out(temp[21]) ) ;
  MUX2_1 mux000022( .i0(SHAMT4[22]), .i1(1'b0), .sel(dataB[4]), .out(temp[22]) ) ;
  MUX2_1 mux000023( .i0(SHAMT4[23]), .i1(1'b0), .sel(dataB[4]), .out(temp[23]) ) ;
  MUX2_1 mux000024( .i0(SHAMT4[24]), .i1(1'b0), .sel(dataB[4]), .out(temp[24]) ) ;
  MUX2_1 mux000025( .i0(SHAMT4[25]), .i1(1'b0), .sel(dataB[4]), .out(temp[25]) ) ;
  MUX2_1 mux000026( .i0(SHAMT4[26]), .i1(1'b0), .sel(dataB[4]), .out(temp[26]) ) ;
  MUX2_1 mux000027( .i0(SHAMT4[27]), .i1(1'b0), .sel(dataB[4]), .out(temp[27]) ) ;
  MUX2_1 mux000028( .i0(SHAMT4[28]), .i1(1'b0), .sel(dataB[4]), .out(temp[28]) ) ;
  MUX2_1 mux000029( .i0(SHAMT4[29]), .i1(1'b0), .sel(dataB[4]), .out(temp[29]) ) ;
  MUX2_1 mux000030( .i0(SHAMT4[30]), .i1(1'b0), .sel(dataB[4]), .out(temp[30]) ) ;
  MUX2_1 mux000031( .i0(SHAMT4[31]), .i1(1'b0), .sel(dataB[4]), .out(temp[31]) ) ;
	
	assign dataOut = (reset)? 32'b0: temp;
	
endmodule