//-----------------------------------------------------------------------------
// Title         : 4-1 multiplexer
//-----------------------------------------------------------------------------

module mux4_32bit( i0, i1, i2, i3, sel, out );
  
  input[31:0] i0, i1, i2, i3 ;
  input[1:0] sel ;
  output[31:0] out ;
  
  assign out = (sel[1])?(sel[0]?i3:i2):(sel[0]?i1:i0) ;
  
endmodule